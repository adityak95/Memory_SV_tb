`include "memory.v"
`include "mem_common.sv"
`include "mem_intf.sv"
`include "mem_tx.sv"
`include "mem_gen.sv"
`include "mem_bfm.sv"
`include "mem_mon.sv"
`include "mem_cov.sv"
`include "mem_sbd.sv"
`include "mem_agent.sv"
`include "mem_env.sv"
`include "mem_assert.sv"
`include "top.sv"
